/* ͬ�� FIFO 4*128  */

// һ��4bit 128��ȵ� ͬ��FIFO���
// @`13
// 2017��6��6��
// ��������ҵ��ѧ�������� EDA�γ����

module fifo(clock,reset,read,write,fifo_in,fifo_out,fifo_empty,fifo_full);

    parameter DEPTH = 128;  						// 128 ��
	 parameter DEPTH_BINARY = 7;  				// ��ȵĶ�����λ��
	 parameter WIDTH = 4;							// 4bit��
	 parameter MAX_CONT = 7'b1111111;			// ���������ֵ127 [0~127]
	 
	 // LED �ƵĶ����Ʊ�ʾ
	 parameter 
		 reg0=7'b0000001,
		 reg1=7'b1001111,
		 reg2=7'b0010010,
		 reg3=7'b0000110,
		 reg4=7'b1001100,
		 reg5=7'b0100100,
		 reg6=7'b0100000,
		 reg7=7'b0001101,
		 reg8=7'b0000000,
		 reg9=7'b0000100,
		 rega=7'b0001000,
		 regb=7'b1100000,
		 regc=7'b0110001,
		 regd=7'b1000010,
		 rege=7'b0110000,
		 regf=7'b0111000;
	 
	 
    input clock,reset,read,write;       			// ʱ�ӣ����ã������أ�д����
    input [WIDTH-1:0]fifo_in;    					// FIFO �������� 
    output[WIDTH-1:0]fifo_out;            	   // FIFO �������
    output fifo_empty,fifo_full;        			// �ձ�־,����־

    reg [WIDTH-1:0]fifo_out;                    // ��������Ĵ���
    reg [WIDTH-1:0]ram[DEPTH-1:0];              // 128��� 8��ȵ� RAM �Ĵ���
    reg [DEPTH_BINARY-1:0]read_ptr,write_ptr,counter;        // ��ָ�룬дָ�룬������ ����Ϊ2^7

    wire fifo_empty,fifo_full;          			// �ձ�־,����־
	 
	 initial                                                
	 begin             
		counter = 0;
		read_ptr = 0;
		write_ptr = 0;
		fifo_out = 0;
	 end              
	 
	 assign fifo_empty = (counter == 0);    		//��־λ��ֵ 
    assign fifo_full = (counter == DEPTH-1);
    
	 always@(posedge clock)    						// ʱ��ͬ������
        if(reset)   										// Reset ����FIFO
            begin
                read_ptr = 0; 
                write_ptr = 0;
                counter = 0;
                fifo_out = 0;                    
            end
        else
            case({read,write})  // ��Ӧ��д����
            2'b00:;  //û�ж�дָ��     
            2'b01:  //дָ���������FIFO                           
            begin
					 if (counter < DEPTH - 1)	// �ж��Ƿ��д
						 begin
						 ram[write_ptr] = fifo_in;
						 counter = counter + 1;
						 write_ptr = (write_ptr == DEPTH-1)?0:write_ptr + 1;
						 end
            end
            2'b10: //��ָ����ݶ���FIFO
            begin
					 if (counter > 0)	// �ж��Ƿ�ɶ�
						 begin
						 fifo_out = ram[read_ptr];
						 counter = counter - 1;
						 read_ptr = (read_ptr == DEPTH-1)?0:read_ptr + 1;
						 end
						 
            end
            2'b11: //��дָ��ͬʱ�����ݿ���ֱ�����
            begin
                if(counter == 0)
                    fifo_out = fifo_in;	// ֱ�����
                else
                begin
                    ram[write_ptr]=fifo_in;
                    fifo_out=ram[read_ptr];
                    write_ptr=(write_ptr==DEPTH-1)?0:write_ptr+1;
                    read_ptr=(read_ptr==DEPTH-1)?0:write_ptr+1;
                end
            end
        endcase
        
endmodule

//module debouncing(
//BJ_CLK,         //�ɼ�ʱ�ӣ�40Hz
//RESET,          //ϵͳ��λ�źŵ͵�ƽ��Ч
//BUTTON_IN,      //���������ź�
//BUTTON_OUT      //�����������ź�
//);
//
//    input BJ_CLK;
//    input RESET;
//    input BUTTON_IN;
//    
//    output BUTTON_OUT;
//
//    reg BUTTON_IN_Q, BUTTON_IN_2Q, BUTTON_IN_3Q;
//    always @(posedge BJ_CLK or negedge RESET)
//    begin
//        if(~RESET)
//            begin
//            BUTTON_IN_Q <= 1'b1;
//            BUTTON_IN_2Q <= 1'b1;
//            BUTTON_IN_3Q <= 1'b1;
//            end
//        else
//            begin   
//            BUTTON_IN_Q <= BUTTON_IN;
//            BUTTON_IN_2Q <= BUTTON_IN_Q;
//            BUTTON_IN_3Q <= BUTTON_IN_2Q;
//            end
//    end
//
//    wire BUTTON_OUT = BUTTON_IN_2Q | BUTTON_IN_3Q;
//
//endmodule
